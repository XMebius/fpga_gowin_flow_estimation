parameter M=8;
parameter N=8;
parameter LATENCY=2;
