`define MODULE_NAME Integer_Division_Top
`define UNSIGNED
`define HAS_REMAINDER
